-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Wed Oct 29 17:02:10 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Maquina_de_estado_secuencia_de_luces IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        A : OUT STD_LOGIC;
        B : OUT STD_LOGIC;
        C : OUT STD_LOGIC;
        D : OUT STD_LOGIC
    );
END Maquina_de_estado_secuencia_de_luces;

ARCHITECTURE BEHAVIOR OF Maquina_de_estado_secuencia_de_luces IS
    TYPE type_fstate IS (S6,S15,S0,S9,S14,S12,S8);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= S0;
            A <= '0';
            B <= '0';
            C <= '0';
            D <= '0';
        ELSE
            A <= '0';
            B <= '0';
            C <= '0';
            D <= '0';
            CASE fstate IS
                WHEN S6 =>
                    reg_fstate <= S15;

                    C <= '1';

                    D <= '0';

                    A <= '0';

                    B <= '1';
                WHEN S15 =>
                    IF ((x = '0')) THEN
                        reg_fstate <= S9;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= S14;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S15;
                    END IF;

                    C <= '1';

                    D <= '1';

                    A <= '1';

                    B <= '1';
                WHEN S0 =>
                    IF ((x = '0')) THEN
                        reg_fstate <= S6;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= S8;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S0;
                    END IF;

                    C <= '0';

                    D <= '0';

                    A <= '0';

                    B <= '0';
                WHEN S9 =>
                    reg_fstate <= S0;

                    C <= '0';

                    D <= '1';

                    A <= '1';

                    B <= '0';
                WHEN S14 =>
                    reg_fstate <= S0;

                    C <= '1';

                    D <= '0';

                    A <= '1';

                    B <= '1';
                WHEN S12 =>
                    IF ((x = '0')) THEN
                        reg_fstate <= S15;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= S14;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S12;
                    END IF;

                    C <= '0';

                    D <= '0';

                    A <= '1';

                    B <= '1';
                WHEN S8 =>
                    reg_fstate <= S12;

                    C <= '0';

                    D <= '0';

                    A <= '1';

                    B <= '0';
                WHEN OTHERS => 
                    A <= 'X';
                    B <= 'X';
                    C <= 'X';
                    D <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
