registro7_inst : registro7 PORT MAP (
		clock	 => clock_sig,
		shiftin	 => shiftin_sig,
		q	 => q_sig
	);
