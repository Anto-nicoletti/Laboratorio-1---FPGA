contador_8_inst : contador_8 PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
