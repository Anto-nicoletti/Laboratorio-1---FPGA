-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Fri Oct 31 18:48:15 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Multiplicador_con_signo IS 
	PORT
	(
		A0 :  IN  STD_LOGIC;
		B0 :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		A1 :  IN  STD_LOGIC;
		CLK :  IN  STD_LOGIC;
		P0 :  OUT  STD_LOGIC;
		P1 :  OUT  STD_LOGIC;
		P2 :  OUT  STD_LOGIC;
		P3 :  OUT  STD_LOGIC;
		NC :  OUT  STD_LOGIC
	);
END Multiplicador_con_signo;

ARCHITECTURE bdf_type OF Multiplicador_con_signo IS 

COMPONENT sumador
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 Cin : IN STD_LOGIC;
		 S : OUT STD_LOGIC;
		 Cout : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_2 <= '0';
SYNTHESIZED_WIRE_37 <= '1';
SYNTHESIZED_WIRE_38 <= '1';



SYNTHESIZED_WIRE_21 <= SYNTHESIZED_WIRE_32 AND SYNTHESIZED_WIRE_33;


b2v_13 : sumador
PORT MAP(A => SYNTHESIZED_WIRE_0,
		 B => SYNTHESIZED_WIRE_34,
		 Cin => SYNTHESIZED_WIRE_2,
		 S => SYNTHESIZED_WIRE_30,
		 Cout => SYNTHESIZED_WIRE_16);


SYNTHESIZED_WIRE_34 <= SYNTHESIZED_WIRE_32 AND SYNTHESIZED_WIRE_35;


SYNTHESIZED_WIRE_14 <= SYNTHESIZED_WIRE_36 AND SYNTHESIZED_WIRE_3;


SYNTHESIZED_WIRE_0 <= SYNTHESIZED_WIRE_36 AND SYNTHESIZED_WIRE_33;


SYNTHESIZED_WIRE_17 <= SYNTHESIZED_WIRE_36 AND SYNTHESIZED_WIRE_4;


SYNTHESIZED_WIRE_4 <= SYNTHESIZED_WIRE_33 AND SYNTHESIZED_WIRE_5;


SYNTHESIZED_WIRE_5 <= NOT(SYNTHESIZED_WIRE_35);



PROCESS(CLK,SYNTHESIZED_WIRE_37,SYNTHESIZED_WIRE_37)
BEGIN
IF (SYNTHESIZED_WIRE_37 = '0') THEN
	SYNTHESIZED_WIRE_35 <= '0';
ELSIF (SYNTHESIZED_WIRE_37 = '0') THEN
	SYNTHESIZED_WIRE_35 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_35 <= A1;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_37,SYNTHESIZED_WIRE_37)
BEGIN
IF (SYNTHESIZED_WIRE_37 = '0') THEN
	SYNTHESIZED_WIRE_32 <= '0';
ELSIF (SYNTHESIZED_WIRE_37 = '0') THEN
	SYNTHESIZED_WIRE_32 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_32 <= B0;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_37,SYNTHESIZED_WIRE_37)
BEGIN
IF (SYNTHESIZED_WIRE_37 = '0') THEN
	SYNTHESIZED_WIRE_33 <= '0';
ELSIF (SYNTHESIZED_WIRE_37 = '0') THEN
	SYNTHESIZED_WIRE_33 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_33 <= A0;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_37,SYNTHESIZED_WIRE_37)
BEGIN
IF (SYNTHESIZED_WIRE_37 = '0') THEN
	SYNTHESIZED_WIRE_36 <= '0';
ELSIF (SYNTHESIZED_WIRE_37 = '0') THEN
	SYNTHESIZED_WIRE_36 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_36 <= B1;
END IF;
END PROCESS;


b2v_inst14 : sumador
PORT MAP(A => SYNTHESIZED_WIRE_14,
		 B => SYNTHESIZED_WIRE_34,
		 Cin => SYNTHESIZED_WIRE_16,
		 S => SYNTHESIZED_WIRE_27,
		 Cout => SYNTHESIZED_WIRE_19);


b2v_inst15 : sumador
PORT MAP(A => SYNTHESIZED_WIRE_17,
		 B => SYNTHESIZED_WIRE_34,
		 Cin => SYNTHESIZED_WIRE_19,
		 S => SYNTHESIZED_WIRE_24,
		 Cout => NC);




SYNTHESIZED_WIRE_3 <= SYNTHESIZED_WIRE_35 XOR SYNTHESIZED_WIRE_33;



PROCESS(CLK,SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_38)
BEGIN
IF (SYNTHESIZED_WIRE_38 = '0') THEN
	P0 <= '0';
ELSIF (SYNTHESIZED_WIRE_38 = '0') THEN
	P0 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	P0 <= SYNTHESIZED_WIRE_21;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_38)
BEGIN
IF (SYNTHESIZED_WIRE_38 = '0') THEN
	P3 <= '0';
ELSIF (SYNTHESIZED_WIRE_38 = '0') THEN
	P3 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	P3 <= SYNTHESIZED_WIRE_24;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_38)
BEGIN
IF (SYNTHESIZED_WIRE_38 = '0') THEN
	P2 <= '0';
ELSIF (SYNTHESIZED_WIRE_38 = '0') THEN
	P2 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	P2 <= SYNTHESIZED_WIRE_27;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_38,SYNTHESIZED_WIRE_38)
BEGIN
IF (SYNTHESIZED_WIRE_38 = '0') THEN
	P1 <= '0';
ELSIF (SYNTHESIZED_WIRE_38 = '0') THEN
	P1 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	P1 <= SYNTHESIZED_WIRE_30;
END IF;
END PROCESS;


END bdf_type;