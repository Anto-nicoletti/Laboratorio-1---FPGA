contador8_inst : contador8 PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
