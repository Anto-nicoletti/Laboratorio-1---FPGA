library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity Multiplicadorbench is
end Multiplicadorbench;

architecture test of Multiplicadorbench is
    signal A0, A1, B0, B1 : std_logic := '0';
    signal P0, P1, P2, P3 : std_logic;

begin

    Suut: entity work.MultiplicadorBlock2
        port map (
            A0 => A0,
            A1 => A1,
            B0 => B0,
            B1 => B1,
            P0 => P0,
            P1 => P1,
            P2 => P2,
            P3 => P3
        );

    -- Proceso de estimulación
    stim_proc: process
    begin
        -- Caso 1: 00 * 00 = 0000
        A1 <= '0'; A0 <= '0';
        B1 <= '0'; B0 <= '0';
        wait for 10 ns;

        -- Caso 2: 01 * 01 = 0001
        A1 <= '0'; A0 <= '1';
        B1 <= '0'; B0 <= '1';
        wait for 10 ns;

        -- Caso 3: 10 * 01 = 0010
        A1 <= '1'; A0 <= '0';
        B1 <= '0'; B0 <= '1';
        wait for 10 ns;

        -- Caso 4: 10 * 10 = 0100
        A1 <= '1'; A0 <= '0';
        B1 <= '1'; B0 <= '0';
        wait for 10 ns;

        -- Caso 5: 11 * 11 = 1001
        A1 <= '1'; A0 <= '1';
        B1 <= '1'; B0 <= '1';
        wait for 10 ns;

        wait; 
    end process;
end test;

