library verilog;
use verilog.vl_types.all;
entity MultiplicadorBlock_vlg_vec_tst is
end MultiplicadorBlock_vlg_vec_tst;
