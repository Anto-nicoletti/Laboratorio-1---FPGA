contador7_inst : contador7 PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
