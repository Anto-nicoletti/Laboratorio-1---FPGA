Library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Sumador is
	port( A : in std_logic;
			B : in std_logic;
			Cin : in std_logic;
			S : out std_logic;
			Cout : out std_logic);
	end Sumador;

architecture comportamiento of Sumador is
		signal sig1: std_logic;
begin
	sig1 <= B xor Cin;
	S <= A XOR sig1;
	COUT <= (A AND Cin) OR (A and B) OR (Cin and B);
end comportamiento;
