contador7_inst : contador7 PORT MAP (
		clock	 => clock_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
