-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Thu Oct 30 20:03:58 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY I2C_maquina_estado IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        sda : IN STD_LOGIC := '0';
        fin_dir : IN STD_LOGIC := '0';
        soy : IN STD_LOGIC := '0';
        fin_dato : IN STD_LOGIC := '0';
        ack : OUT STD_LOGIC;
        hab_dir : OUT STD_LOGIC;
        hab_dat : OUT STD_LOGIC
    );
END I2C_maquina_estado;

ARCHITECTURE BEHAVIOR OF I2C_maquina_estado IS
    TYPE type_fstate IS (Oscioso,Guardar_dir,R_W,AC,guardar_dato);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,sda,fin_dir,soy,fin_dato)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Oscioso;
            ack <= '0';
            hab_dir <= '0';
            hab_dat <= '0';
        ELSE
            ack <= '0';
            hab_dir <= '0';
            hab_dat <= '0';
            CASE fstate IS
                WHEN Oscioso =>
                    IF ((sda = '1')) THEN
                        reg_fstate <= Oscioso;
                    ELSIF ((sda = '0')) THEN
                        reg_fstate <= Guardar_dir;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Oscioso;
                    END IF;

                    hab_dat <= '0';

                    hab_dir <= '0';

                    ack <= '0';
                WHEN Guardar_dir =>
                    IF (((fin_dir = '1') AND (soy = '0'))) THEN
                        reg_fstate <= Oscioso;
                    ELSIF ((fin_dir = '0')) THEN
                        reg_fstate <= Guardar_dir;
                    ELSIF (((fin_dir = '1') AND (soy = '1'))) THEN
                        reg_fstate <= R_W;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guardar_dir;
                    END IF;

                    hab_dat <= '0';

                    hab_dir <= '1';

                    ack <= '0';
                WHEN R_W =>
                    reg_fstate <= AC;

                    hab_dat <= '0';

                    hab_dir <= '0';

                    ack <= '0';
                WHEN AC =>
                    reg_fstate <= guardar_dato;

                    hab_dat <= '0';

                    hab_dir <= '0';

                    ack <= '1';
                WHEN guardar_dato =>
                    IF ((fin_dato = '0')) THEN
                        reg_fstate <= guardar_dato;
                    ELSIF ((fin_dato = '1')) THEN
                        reg_fstate <= Oscioso;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= guardar_dato;
                    END IF;

                    hab_dat <= '1';

                    hab_dir <= '0';

                    ack <= '0';
                WHEN OTHERS => 
                    ack <= 'X';
                    hab_dir <= 'X';
                    hab_dat <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
