library verilog;
use verilog.vl_types.all;
entity Multiplicador_con_signo_Block_vlg_check_tst is
    port(
        NC              : in     vl_logic;
        P0              : in     vl_logic;
        P1              : in     vl_logic;
        P2              : in     vl_logic;
        P3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Multiplicador_con_signo_Block_vlg_check_tst;
