registro8_inst : registro8 PORT MAP (
		clock	 => clock_sig,
		shiftin	 => shiftin_sig,
		q	 => q_sig
	);
