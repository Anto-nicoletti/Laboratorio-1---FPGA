library verilog;
use verilog.vl_types.all;
entity opcion_multi_vlg_vec_tst is
end opcion_multi_vlg_vec_tst;
