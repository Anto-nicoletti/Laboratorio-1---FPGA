contador_8_inst : contador_8 PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
