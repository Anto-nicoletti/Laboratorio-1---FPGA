library verilog;
use verilog.vl_types.all;
entity SumadorBlock1_vlg_vec_tst is
end SumadorBlock1_vlg_vec_tst;
